module AG(input  [31:0] SrcAE, SrcBE,output [31:0] AGOut);
	assign AGOut = SrcAE + SrcBE;
endmodule